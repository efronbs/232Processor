`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Rose-Hulman CSSE dept. (student)
// Engineer: Thomas Bonatti
// 
// Create Date:    01/28/2015 
// Design Name: 
// Module Name:    ALU16bit 
// Project Name: 	csse232 comp arc final project (team B)
//
//
//////////////////////////////////////////////////////////////////////////////////
module mainRegAdrs(adrsOut
    );
	output reg [2:0] adrsOut = 0;

endmodule
