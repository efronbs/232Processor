`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Rose-Hulman CSSE dept. (student)
// Engineer: Thomas Bonatti
// 
// Create Date:    01/28/2015 
// Design Name: 
// Module Name:    ALU16bit 
// Project Name: 	csse232 comp arc final project (team B)
//
//
//////////////////////////////////////////////////////////////////////////////////
module adder16bit(aIn, bIn, outPin
    );
	input [15:0] aIn, bIn;
	output reg [15:0] outPin;

	always @(aIn, bIn) begin
		outPin = aIn + bIn;
	end

endmodule
